/*
This module contains our processor that calculates important signals for our game
*/
`include "pc4/skeleton.v"
module processingUnit(clock, reset);
	input clock, reset;
//	output [4:0] ctrl_writeReg;
//	output ctrl_writeEnable;
//	output [31:0] data_writeReg;
	
	skeleton my_processor(.clock(clock), .reset(reset)); 
	//outputs will be changed	
		
		
		
		
		
		
		
endmodule