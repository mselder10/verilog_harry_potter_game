module letter(letter, clk, row, col,
			  get_ready, times_up, leaderboard);
	
	input clk, get_ready, times_up, leaderboard;
	input [8:0] row;
	input [9:0] col;

	wire [4:0] get_ready_letter, times_up_letter, house_cup_letter;
	wire [4:0] display_letter;

	wire [4:0] get_ready_ADDR, times_up_ADDR, house_cup_ADDR;
	wire [12:0] ADDR;
	wire [15:0] offset_ADDR;

	output letter;

	// get ready logic
	get_ready 	readyz(.row(row), .col(col), .clk(clk),
					   .letter(get_ready_letter), .pixel(get_ready_ADDR));

	time_is_up 	timez(.row(row), .col(col), .clk(clk), 
					  .letter(times_up_letter), .pixel(times_up_ADDR));

	house_cup 	cupz( .row(row), .col(col), .clk(clk), .leaderboard(leaderboard),
				   	  .letter(house_cup_letter), .pixel(house_cup_ADDR));

	// what to display
	assign display_letter = get_ready 	 ? get_ready_letter : 5'dz;
	assign display_letter = times_up  	 ? times_up_letter  : 5'dz;
	assign display_letter = leaderboard  ? house_cup_letter : 5'dz;

	assign ADDR = get_ready 	 ? get_ready_ADDR : 12'dz;
	assign ADDR = times_up  	 ? times_up_ADDR  : 12'dz;
	assign ADDR = leaderboard  	 ? house_cup_ADDR : 12'dz;

	// find letter offset in mif file
	assign offset_ADDR = ADDR + display_letter*2500;

	letters alphabet(.address(offset_ADDR),
				   	 .clock(~clk),
				   	 .q(letter));

endmodule