module trace_change(trace_to_display, clk, p1_traced, p2_traced, trace_screen_on, end_game_early, trace_count, previous_trace_displayed, two_player_mode);
	
	input trace_screen_on, clk, two_player_mode;
	input [15:0] p1_traced, p2_traced;
	
	output reg [5:0] trace_count;
	reg [15:0] trace0, trace1, trace2, trace3, trace4;
	
	output reg [15:0] trace_to_display, previous_trace_displayed;
	output reg end_game_early;
	
	initial begin
		trace_count <= 0;
		trace_to_display <= 16'h0231;
		end_game_early <= 0;
		trace1 <= 16'h0075;
		trace2 <= 16'h8ca9;	
		trace3 <= 16'h8f23;
		trace4 <= 16'hd9be;
	end
	
	always@(posedge clk & trace_screen_on)
	begin
		// if user trace and trace display are the same, change the trace displayed
		if((p1_traced & trace_to_display)==trace_to_display || (((p2_traced & trace_to_display)==trace_to_display) & two_player_mode))
		begin
			trace_count = trace_count + 1;
			if(trace_count == 1)
			begin
				//previous_trace_displayed <= trace_to_display;
				trace_to_display <= trace1;
			end
			else if (trace_count == 2)
			begin
				//previous_trace_displayed <= trace_to_display;
				trace_to_display <= trace2;
			end
			else if (trace_count == 3)
			begin
				//previous_trace_displayed <= trace_to_display;
				trace_to_display <= trace3;
			end
			else if (trace_count == 4)
			begin
				//previous_trace_displayed <= trace_to_display;
				trace_to_display <= trace4;
			end
			else if (trace_count == 5)
			begin
				trace_count <= 0;
				end_game_early <= 1;
			end
		end
		
	end

endmodule 